
module eced4260beamformer(


);










endmodule







