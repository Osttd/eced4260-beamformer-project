

module delaybeamerformer_tb();









endmodule












